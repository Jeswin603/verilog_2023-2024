library verilog;
use verilog.vl_types.all;
entity jhonson_counter_tb is
end jhonson_counter_tb;
