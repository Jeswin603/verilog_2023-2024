library verilog;
use verilog.vl_types.all;
entity decodertwo_tb is
end decodertwo_tb;
