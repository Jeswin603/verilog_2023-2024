library verilog;
use verilog.vl_types.all;
entity dexfour_tb is
end dexfour_tb;
