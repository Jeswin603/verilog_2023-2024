library verilog;
use verilog.vl_types.all;
entity dfliptb is
end dfliptb;
