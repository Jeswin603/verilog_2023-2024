library verilog;
use verilog.vl_types.all;
entity free_runner_tb is
end free_runner_tb;
