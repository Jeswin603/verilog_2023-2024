module anand(
input a,b,
output c);
assign y =~(a&b);
endmodule
