module not1(
input a,
output c );
assign c = ~a;
endmodule


