library verilog;
use verilog.vl_types.all;
entity twomux_tb is
end twomux_tb;
