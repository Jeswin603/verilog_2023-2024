library verilog;
use verilog.vl_types.all;
entity demuxtwo_tb is
end demuxtwo_tb;
