library verilog;
use verilog.vl_types.all;
entity twomuxtb is
end twomuxtb;
