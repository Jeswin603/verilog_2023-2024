library verilog;
use verilog.vl_types.all;
entity not1 is
    port(
        a               : in     vl_logic;
        c               : out    vl_logic
    );
end not1;
